library verilog;
use verilog.vl_types.all;
entity proj3342_vlg_vec_tst is
end proj3342_vlg_vec_tst;
